module muxValor(
    input v1, v0, 
    output [12:0] valor
    );

endmodule