module adder_sub_12bit(
    input [11:0] a, b, cin,
    output [11:0] sum, cout
);

    wire carry[12:0];
    assign

    genvar i;
    generate 
        for (i = 0, i<12, i = i+ 1) begin adder_chain 

        end

    endgenerate

endmodule