module registerD12bit(
    input clk, rst, d_ld, d_clr,
    input [11:0] d_in,
    output reg [11:0] q);

    always@(posedge clk or posedge rst) begin 
        
    end
endmodule