module piscaled(input clk, c);

endmodule