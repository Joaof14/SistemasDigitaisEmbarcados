module datapath(
    input clk, rst,

    //entradas do datapath

    //entradas de sinais de comando

    //saídas de sinais de status

    //saídas de dados
)