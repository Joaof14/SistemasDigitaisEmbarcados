module comparators(
    input [11:0] d, 
    output m
);
    

endmodule