module control_unit(
    input clk, rst
    //entradas de controle

    //sinais de status

    //sinais de comando

    //saida de controle
);

endmodule