module adder_sub_1bit(
    input a, b, cin,
    output sum, cout
);

endmodule