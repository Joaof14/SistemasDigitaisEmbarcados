module muxValorMoeda(
    input S, s0, s1, 
    output [12:0] valor
    );
endmodule