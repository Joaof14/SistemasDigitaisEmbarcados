module comparators();

endmodule